.title KiCad schematic
L4 Net-_C4-Pad1_ Net-_C5-Pad1_ 200n
L3 Net-_C3-Pad1_ Net-_C4-Pad1_ 200n
C4 Net-_C4-Pad1_ GND 67p
L5 Net-_C5-Pad1_ /sig_out 200n
C5 Net-_C5-Pad1_ GND 67p
J2 /sig_out GND Conn_Coaxial
C6 /sig_out GND 67p
R2 /sig_out GND 50R
C3 Net-_C3-Pad1_ GND 67p
C1 Net-_C1-Pad1_ GND 67p
J1 /sig_in GND Conn_Coaxial
R1 /sig_in Net-_C1-Pad1_ 50R
L1 Net-_C1-Pad1_ Net-_C2-Pad1_ 200n
C2 Net-_C2-Pad1_ GND 67p
L2 Net-_C2-Pad1_ Net-_C3-Pad1_ 200n
.end
