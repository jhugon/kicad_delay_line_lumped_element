.title KiCad schematic
J1 /sig_in GND Conn_Coaxial
L4 Net-_C4-Pad1_ Net-_C5-Pad1_ 200n
L3 Net-_C3-Pad1_ Net-_C4-Pad1_ 200n
C4 Net-_C4-Pad1_ unconnected-_C4-Pad2_ 67p
C1 /sig_in unconnected-_C1-Pad2_ 67p
L5 Net-_C5-Pad1_ /sig_out 200n
L1 /sig_in Net-_C2-Pad1_ 200n
C2 Net-_C2-Pad1_ unconnected-_C2-Pad2_ 67p
L2 Net-_C2-Pad1_ Net-_C3-Pad1_ 200n
C3 Net-_C3-Pad1_ unconnected-_C3-Pad2_ 67p
C5 Net-_C5-Pad1_ unconnected-_C5-Pad2_ 67p
C6 /sig_out unconnected-_C6-Pad2_ 67p
J2 /sig_out GND Conn_Coaxial
.end
